* ============================================================================
* SKY130 Multi-Vth Device Models for Ternary Logic - TT Corner
* ============================================================================
* GT-LOGIC Ternary CMOS Cell Library
* Extracted from SkyWater SKY130 Open PDK
* Corner: Typical-Typical (TT) @ 30C nominal
* ============================================================================

* MISMATCH PARAMETERS (all set to 0 for TT corner)
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_slope = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_slope = 0.0

.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__nfactor_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__toxe_slope = 0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope = 0.0
.param sky130_fd_pr__nfet_01v8__voff_slope = 0.0
.param sky130_fd_pr__nfet_01v8__nfactor_slope = 0.0

.param sky130_fd_pr__pfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__toxe_slope = 0.0
.param sky130_fd_pr__pfet_01v8__vth0_slope = 0.0
.param sky130_fd_pr__pfet_01v8__voff_slope = 0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope = 0.0

.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope = 0.0

* DEVICE MODELS (BSIM4)
.include "E:/Tritone-V2/tritone-complete/pdk/sky130_fd_pr/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.pm3.spice"
.include "E:/Tritone-V2/tritone-complete/pdk/sky130_fd_pr/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.pm3.spice"
.include "E:/Tritone-V2/tritone-complete/pdk/sky130_fd_pr/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.pm3.spice"
.include "E:/Tritone-V2/tritone-complete/pdk/sky130_fd_pr/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.pm3.spice"
