* ============================================================================
* MULTI-CORNER BSIM4 PVT CHARACTERIZATION - Multi-Vth STI for SKY130
* ============================================================================
* GT-LOGIC Ternary CMOS Cell Library
*
* Sweeps all 5 process corners (TT, SS, FF, SF, FS) with voltage and
* temperature variations for complete PVT characterization.
*
* Run in Docker: ngspice -b tb_sti_multicorner_bsim4.spice
* ============================================================================

* ============================================================================
* CONTROL SCRIPT FOR MULTI-CORNER ANALYSIS
* ============================================================================
.control

set filetype = ascii
set wr_vecnames

echo "================================================================"
echo "SKY130 BSIM4 Multi-Corner STI Characterization"
echo "================================================================"
echo ""
echo "Process Corners: TT, SS, FF, SF, FS"
echo "Voltage Range: 1.62V to 1.98V (1.8V ±10%)"
echo "Temperature Range: -40C to 125C"
echo ""

* Create results directory
shell mkdir -p /tritone/spice/results

* ============================================================================
* Define corner simulation function
* ============================================================================

* We'll run each corner as a separate netlist since ngspice
* doesn't support dynamic model switching well

* First, generate individual corner testbenches
foreach corner tt ss ff sf fs

  echo ""
  echo "================================================================"
  echo "Processing $corner corner..."
  echo "================================================================"

  * Create corner-specific netlist
  shell cat > /tritone/spice/results/run_$corner.spice << CORNER_EOF
* SKY130 Multi-Vth STI - $corner Corner
* Auto-generated multi-corner testbench

* Include SKY130 BSIM4 models
.include "/tritone/pdk/sky130_fd_pr/models/corners/$corner.spice"

* Include the redesigned STI cell
.include "/tritone/spice/cells/sti_multivth_sky130.spice"

* Power supplies
VVDD vdd 0 DC 1.8
VVSS vss 0 DC 0

* Input
VIN in 0 DC 0

* DUT
XDUT in out vdd vss STI_MULTIVTH_SKY130

* Load
CL out 0 10f

.control
set filetype = ascii

echo "=== $corner Corner @ 27C, VDD=1.8V ==="

* DC sweep
dc VIN 0 1.8 0.005

* Save data
wrdata /tritone/spice/results/dc_$corner.dat v(out)

* Key measurements
meas dc vout_low FIND v(out) AT=0
meas dc vout_mid FIND v(out) AT=0.9
meas dc vout_high FIND v(out) AT=1.8
meas dc vil_th WHEN v(out)=1.35 CROSS=1
meas dc vih_th WHEN v(out)=0.45 CROSS=1

let vmid_err = abs(vout_mid - 0.9)
let nml = vil_th
let nmh = 1.8 - vih_th

echo "Results:"
echo "  Vout(0V)=$&vout_low Vout(0.9V)=$&vout_mid Vout(1.8V)=$&vout_high"
echo "  VIL=$&vil_th VIH=$&vih_th"
echo "  Mid-error=$&vmid_err NML=$&nml NMH=$&nmh"

* Temperature variations
echo ""
echo "--- Temperature Sweep ---"

set temp = -40
dc VIN 0 1.8 0.01
meas dc vmid_m40 FIND v(out) AT=0.9
let err_m40 = abs(vmid_m40 - 0.9)
echo "  -40C: Vmid=$&vmid_m40 err=$&err_m40"

set temp = 85
dc VIN 0 1.8 0.01
meas dc vmid_85 FIND v(out) AT=0.9
let err_85 = abs(vmid_85 - 0.9)
echo "   85C: Vmid=$&vmid_85 err=$&err_85"

set temp = 125
dc VIN 0 1.8 0.01
meas dc vmid_125 FIND v(out) AT=0.9
let err_125 = abs(vmid_125 - 0.9)
echo "  125C: Vmid=$&vmid_125 err=$&err_125"

set temp = 27

* Voltage variations
echo ""
echo "--- Voltage Sweep ---"

alter VVDD = 1.62
dc VIN 0 1.62 0.01
meas dc vmid_lv FIND v(out) AT=0.81
let err_lv = abs(vmid_lv - 0.81)
echo "  VDD=1.62V: Vmid=$&vmid_lv err=$&err_lv"

alter VVDD = 1.98
dc VIN 0 1.98 0.01
meas dc vmid_hv FIND v(out) AT=0.99
let err_hv = abs(vmid_hv - 0.99)
echo "  VDD=1.98V: Vmid=$&vmid_hv err=$&err_hv"

quit
.endc
.end
CORNER_EOF

  * Run the corner simulation
  shell ngspice -b /tritone/spice/results/run_$corner.spice > /tritone/spice/results/log_$corner.txt 2>&1

  echo "Saved results to /tritone/spice/results/log_$corner.txt"

end

* ============================================================================
* SUMMARY REPORT
* ============================================================================
echo ""
echo "================================================================"
echo "MULTI-CORNER CHARACTERIZATION COMPLETE"
echo "================================================================"
echo ""
echo "Results saved in /tritone/spice/results/"
echo ""
echo "Corner Summary:"

foreach corner tt ss ff sf fs
  echo ""
  echo "--- $corner ---"
  shell grep -A3 "Results:" /tritone/spice/results/log_$corner.txt 2>/dev/null || echo "  (check log file)"
end

echo ""
echo "================================================================"
echo "DATA FILES GENERATED:"
echo "================================================================"
shell ls -la /tritone/spice/results/*.dat 2>/dev/null || echo "  (no .dat files)"
echo ""

quit

.endc

* Dummy circuit (control script runs the actual simulations)
V1 dummy 0 DC 0
R1 dummy 0 1k

.end
